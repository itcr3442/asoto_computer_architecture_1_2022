`ifndef TYPES_SV
`define TYPES_SV

typedef logic[3:0]   nibble;
typedef logic[15:0]  hword;
typedef logic[31:0]  word;
typedef logic[63:0]  dword;
typedef logic[127:0] qword;
typedef logic[30:0]  hptr;
typedef logic[29:0]  ptr;
typedef logic[27:0]  qptr;

`endif
