`include "core/uarch.sv"

module core_alu
#(parameter W=16)
(
	input  logic          clk,
	                      rst_n,

	input  insn_decode    dec,
	input  logic          start,
	input  logic[W - 1:0] a,
	                      b,

	output wb_line        wb,
	output hword          raw_mask
);

	logic[W - 1:0] b_or_imm, q;

	assign b_or_imm = dec.data.uses_imm ? {{(W - 6){dec.data.imm[5]}}, dec.data.imm} : b;

	core_raw_mask rd_mask
	(
		.r(dec.data.rd),
		.enable(start),
		.*
	);

	always_comb
		unique case(dec.alu.op)
			`ALU_AND:
				q = a & b;

			`ALU_ORR:
				q = a | b;

			`ALU_XOR:
				q = a ^ b;

			`ALU_SHL:
				q = a << b_or_imm;

			`ALU_SHR:
				q = a >> b_or_imm;

			`ALU_ADD:
				q = a + b_or_imm;

			`ALU_SUB:
				q = a - b_or_imm;

`ifdef VERILATOR
			0: ;
`endif
		endcase

	always @(posedge clk or negedge rst_n)
		if(!rst_n) begin
			wb <= {$bits(wb_line){1'bx}};
			wb.ready <= 0;
		end else begin
			wb.rd <= dec.data.rd;
			wb.value <= q;
			wb.ready <= start;
		end

endmodule
